[{"type":"Toc","source_relative_path":"obj/api/toc.yml","output":{".html":{"relative_path":"api/toc.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\zr3rjvdp.cwm","hash":"Ue9e8GsRaRMMaJ/7r4I21iwBtxbGCYZ3enprAH/472w="}},"is_incremental":false,"version":""},{"type":"Toc","source_relative_path":"toc.yml","output":{".html":{"relative_path":"toc.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\xv45y5gd.21g","hash":"Oa9PuD4E1hvZnCkVjUgzNBX6S00Zo5YilamTERTZo54="}},"is_incremental":false,"version":""},{"type":"Toc","source_relative_path":"articles/toc.md","output":{".html":{"relative_path":"articles/toc.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\jh1g1usi.pfr","hash":"BlPxk5mtl2kgfcZUgkEguqiSAR/EUyUTT4EdebwkQvs="}},"is_incremental":false,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.CladdingType.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.CladdingType.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\5snt5hyg.vci","hash":"lVS9on7Ko+6wjhxQOYQ/kRsoPmAYDMuUQkM9eYDbxnQ="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.BillboardSide.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.BillboardSide.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\rdvcmdnv.dxf","hash":"AMMx5qKe1gSsBs0c2qufw2/Yz8QoPHkB/4H3MCgcgUQ="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\zwt1kqkg.2yv","hash":"WD6T6dPQLvV65Ao32Jj1jsPUQKQikNcl5XS6HaG40Rs="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"index.md","output":{".html":{"relative_path":"index.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\rfhhyqkf.cfz","hash":"GGOovSab6ZFxRkwbTiKX/AxcXz9WU1qSZOSIhjRqq74="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"api/index.md","output":{".html":{"relative_path":"api/index.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\kfgkzdvw.zap","hash":"ZcRFJgNhvhM6kAH28Vkb5TxxGPe7FlftmernEpHWKBw="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.LiftPoint.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.LiftPoint.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\haxnoexw.4kx","hash":"UWuSbbua29M0lCcdJnF13flXgIsnZxwnLbm2cm3NQXc="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Flashing.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Flashing.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\ifa41nep.pqz","hash":"/Z1Yqni1xE1MtVBT8Ig82/yJOtenhBSmqIZ1CjJEmaM="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/BeamApplication.Properties.yml","output":{".html":{"relative_path":"api/BeamApplication.Properties.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\z5idyn1c.z02","hash":"h/nL0cxofZ70zmMRVgrRntGncFFmSh/FcFUb/erqg/0="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.HorizontalRailing.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.HorizontalRailing.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\wpzkvpmq.u5p","hash":"vdMnmvgD7Kgdm1DYydu19eFlO4kGTZROe/kbIVCo7Yw="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.GalHole.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.GalHole.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\y5s5u2hw.vsk","hash":"U52jU16g1qRmFEc2/6Un52l4fRguiTtdmIKoY6V5Z0o="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Frame.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Frame.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\5erx3x4s.dok","hash":"YjqD+jzBBjal9OuF+I0MSAbCdjuSo7dRg+PzsCDwyrw="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"articles/intro.md","output":{".html":{"relative_path":"articles/intro.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\u5mjeks4.eyz","hash":"yF4cM99miGSsrT64oV0kgkl56YkQylthgw5Gl1aJqzo="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.BetterEASupport.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.BetterEASupport.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\cxiwoky0.u21","hash":"o8N4ToU3YK3vHGCchaPhyaDiWY1y0R8cxwhVzhKZBqY="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid._3DFascia.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid._3DFascia.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\n4mb5wlv.m5l","hash":"CqhrY+n9Zw7NgN1JQ1RatViWPBXHA31FwrO2yQDcgg4="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Walkway.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Walkway.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\qtgps3dk.spf","hash":"3p6YwhRNoU1QNP0VJ3YbUBuri2XQwl4z0Mpspun2XB4="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Hatch.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Hatch.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\se0yoai4.r2l","hash":"aT2gJvABTU/SNV/MqeIW/AFGhJaraTxc919CjB5kYtg="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Cladding.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Cladding.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\dj40phno.s5j","hash":"dVYOcgCzxg3NWvMT0Ns0QgjRvITlQtQTuTlTD6ZXpaU="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Plate.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Plate.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\m0g5pufp.jrb","hash":"p64FLssi3NwAtaYd4AA15zL+25JJpzIPi/e2QgSwOaE="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/BeamApplication.Properties.Resources.yml","output":{".html":{"relative_path":"api/BeamApplication.Properties.Resources.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\vxkmj2th.wd0","hash":"bPB7q08h+JETXPb5QMwhAo/77Hw1pd307iAXbd3gv70="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Colour.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Colour.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\20aqm1ce.bbe","hash":"g/6yjeyWlGXJMMmQVddUHLuX2+V6Eo1WKqXNgfTyv0Y="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Diagonal.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Diagonal.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\quyipvtv.wzy","hash":"k35q6MkBX52DUWw25chmNWuuMBalGqu21mzHI4pGUcI="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.HorizontalBeam.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.HorizontalBeam.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\jlsmt1db.swj","hash":"Q+4hlm5Z6RJ5Lr2dMnu0ylKWPnw28HHeJYttLBH2UHw="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.ModelParameters.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.ModelParameters.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\vwmepu5f.ros","hash":"7Eu7HPtLgfFloeWqX/Zsw305ffBX27bEleZKWkg3osY="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.FasciaBox.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.FasciaBox.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\sbgaj00j.c5h","hash":"9ZK9mvQnfFT6teyxMehkQ3uJ4dgIuWSSM09EzkANYH4="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.ZBracket.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.ZBracket.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\lsowr2iu.1jp","hash":"Ob7r8SEgRDcZ2Z8ceM97Fmx2m2w2gXVNUmnIZPzQxKw="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Waler.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Waler.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\yrpaqkup.evd","hash":"7nbCfGyAKqaEn1PdABQ7Slq7kC7gynp3LbdFUyNZLXI="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.LadderBuilder.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.LadderBuilder.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\q0k24grc.2qp","hash":"drUEiPt4dx3cTx+ojBfTlsNLje9O0Zqz+JRTbV6LRQU="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Box.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Box.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\sg2pcqes.pdl","hash":"cOrPZGbC93ZdssTv8XdRLegM+BvVqp62eC9YwiSIkyA="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.CameraArm.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.CameraArm.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\rduta2px.smd","hash":"Tz9ekHpwVYzw2r6Nw0tSa/jBmEOZJ2Nesorz7Qiod6Y="}},"is_incremental":true,"version":""},{"type":"ManagedReference","source_relative_path":"obj/api/TeklaBillboardAid.Form1.yml","output":{".html":{"relative_path":"api/TeklaBillboardAid.Form1.html","link_to_path":"C:\\Users\\Thomas\\Documents\\Uni\\JFC\\Code\\ALL CODES\\MAIN CODING\\obj\\.cache\\build\\bb0zjbvt.qc3\\s4ebobla.nxj","hash":"nv68PIYSLgELmpwNsvi9gxnZPROEbLb3hQAH0M+5eWg="}},"is_incremental":true,"version":""}]